module main

import levenshtein

fn main(){
	println(levenshtein.calculate("voiture","voilure"))
}